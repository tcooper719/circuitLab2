module AND1 (output oand1, input A, B);
    assign oand1 = A & B;//this assigns the output oand1 to 
endmodule