module NOT1 (output wire onot1, input A);
    assign onot1 = ~A;//this assigns the output A to 
endmodule 