module NOT (output wire onot, input A);
    assign onot = ~A;//this assigns the output A to 
endmodule 